module and_gate (
	input a, b,		// Defining inputs A & B of AND Gate
	output out		// Defining output of AND Gate
);

assign out = a & b;	// Logic Implementation

endmodule
